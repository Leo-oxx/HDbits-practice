//创建一个实现非门的模块。
module top_module( input in, output out );

	assign out = ~in;
	
endmodule