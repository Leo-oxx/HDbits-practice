//创建一个有一个输入和一个输出的模块，其行为类似于导线。
module top_module( input in, output out );
	assign out = in;
endmodule