//建立一个没有输入、只有一个输出且输出恒为 0 的电路
module top_module(output zero);// Module body starts after semicolon
    assign zero = 0;
endmodule
