//给定几个输入向量，将它们连接起来，然后分割成几个输出向量。
//有六个 5 位输入向量：a、b、c、d、e 和 f，总共 30 位输入。
//有四个 8 位输出向量：w、x、y 和 z，共 32 位输出。输出应该是输入向量的连接，后面跟两个 1 位：

module top_module (
    input [4:0] a, b, c, d, e, f,
    output [7:0] w, x, y, z );//

    assign w[7:0] = {a[4:0], b[4:2]};// 5 + 3
	assign x[7:0] = {b[1:0], c[4:0], d[4]};//2 + 5 + 1
	assign y[7:0] = {d[3:0], e[4:1]};//4 + 4
	assign z[7:0] = {e[0], f[4:0], 2'b11};//1 + 5 + 2

endmodule
